`timescale 1ns/100ps

module testbench();

   
endmodule
/*
        ex_MULT_busy_out_tb         == ex_MULT_busy_out &&
        ex_CDB_arb_stall_out_tb     == ex_CDB_arb_stall_out &&
        ex_branch_mispredict_out_tb == ex_branch_mispredict_out &&
        ex_branch_inst_out_tb       == ex_branch_inst_out &&
        ex_store_inst_out_tb        == ex_store_inst_out &&
        ex_CDB_tag_out              == ex_CDB_tag_out &&
        ex_ROB_number_out           == ex_ROB_number_out &&
        ex_result_out_tb            == ex_result_out &&
        ex_NPC_out_tb               == ex_NPC_out */
